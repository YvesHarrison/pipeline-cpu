module get_switch(number,switch);
	input	[4:0]	switch;
	output	[7:0]	number;

	//assign lcd[0]=switch[0];
	//assign lcd[1]=switch[1];
	//assign lcd[2]=switch[2];
	//assign lcd[3]=switch[3];
	//assign lcd[4]=switch[4];
	assign	number[4]=switch[4];
	assign	number[3]=switch[3];
	assign	number[2]=switch[2];
	assign 	number[1]=switch[1];
	assign	number[0]=switch[0];
	
endmodule